module Graphic_EQ (
	CLOCK_50,
	reset,
	AUD_ADCDAT,

	AUD_BCLK,
	AUD_ADCLRCK,
	AUD_DACLRCK,

	AUD_XCK,
	AUD_DACDAT,
	I2C_SCLK,
	I2C_SDAT,
	
	set,
	bass_level,
	mid_level,
	treble_level
);

	input CLOCK_50, reset, AUD_ADCDAT,set;
	inout AUD_BCLK, AUD_ADCLRCK, AUD_DACLRCK,I2C_SCLK,I2C_SDAT;
	output AUD_XCK, AUD_DACDAT;
	
	input signed [4:0] bass_level,mid_level,treble_level;
	
	wire [31:0] l_channel_audio_in, r_channel_audio_in, l_channel_audio_out, r_channel_audio_out;
	wire read_ready, write_ready, read_enable, write_enable;
	wire read_clock;
	wire [9:0] bass_ctrl, low_mid_ctrl, mid_ctrl, treble_ctrl;
	
	assign read_enable = read_ready;
	assign write_enable = write_ready;

	Audio_Controller audioAudio_Controller(
		// Inputs
		.CLOCK_50(CLOCK_50),
		.reset(~reset),

		.read_audio_in(1'b1),
		.left_channel_audio_out(l_channel_audio_out),
		.right_channel_audio_out(r_channel_audio_out),
		.write_audio_out(1'b1),

		.AUD_ADCDAT(AUD_ADCDAT),

		// Bidirectionals
		.AUD_BCLK(AUD_BCLK),
		.AUD_ADCLRCK(AUD_ADCLRCK),
		.AUD_DACLRCK(AUD_DACLRCK),

		// Outputs
		.left_channel_audio_in(l_channel_audio_in),
		.right_channel_audio_in(r_channel_audio_in),
		.audio_in_available(read_ready),

		.audio_out_allowed(write_ready),

		.AUD_XCK(AUD_XCK),
		.AUD_DACDAT(AUD_DACDAT)
	);


	avconf conf(
		//	Host Side
						.CLOCK_50(CLOCK_50),
						.reset(reset),
						//	I2C Side
						.I2C_SCLK(I2C_SCLK),
						.I2C_SDAT(I2C_SDAT)
	);

equalizer_ctrl eq_left(
	.enter(set),
	
	.bass_level(bass_level),
	.mid_level(mid_level),
	.treble_level(treble_level),

	.d_in(l_channel_audio_in),
	.d_out(l_channel_audio_out),
	.clk(read_ready));
	
equalizer_ctrl eq_right(
	.enter(set),
	
	.bass_level(bass_level),
	.mid_level(mid_level),
	.treble_level(treble_level),

	.d_in(r_channel_audio_in),
	.d_out(r_channel_audio_out),
	.clk(read_ready));
	
endmodule
